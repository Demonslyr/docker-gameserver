#
# LinuxGSM Valheim Dockerfile
#
# https://github.com/Demonslyr/docker-gameserver
#

FROM docker.atriarch.systems/linuxgsm:ubuntu-2204
LABEL maintainer="Atriarch Systems <postmaster@mail.atriarch.systems>"
ARG SHORTNAME=vh
ENV GAMESERVER=vhserver

WORKDIR /app

## Auto install game server requirements
RUN depshortname=$(curl --connect-timeout 10 -s https://cdn.atriarch.systems/File/cdn-wfe/ab91225aa4ee457899a9e0368e253ebd |awk -v shortname="vh" -F, '$1==shortname {$1=""; print $0}') \
  && if [ -n "${depshortname}" ]; then \
  echo "**** Install ${depshortname} ****" \
  && apt-get update \
  && apt-get install -y ${depshortname} \
  && apt-get -y autoremove \
  && apt-get clean \
  && rm -rf /var/lib/apt/lists/* /tmp/* /var/tmp/*; \
  fi

HEALTHCHECK --interval=1m --timeout=1m --start-period=2m --retries=1 CMD /app/entrypoint-healthcheck.sh || exit 1

RUN date > /build-time.txt

ENTRYPOINT ["/bin/bash", "./entrypoint.sh"]
